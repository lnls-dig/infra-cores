`define ADDR_AFC_MGMT_CLK_DISTRIB      3'h0
`define AFC_MGMT_CLK_DISTRIB_SI57X_OE_OFFSET 0
`define AFC_MGMT_CLK_DISTRIB_SI57X_OE 32'h00000001
`define AFC_MGMT_CLK_DISTRIB_RESERVED_OFFSET 1
`define AFC_MGMT_CLK_DISTRIB_RESERVED 32'hfffffffe
`define ADDR_AFC_MGMT_DUMMY            3'h4
`define AFC_MGMT_DUMMY_RESERVED_OFFSET 0
`define AFC_MGMT_DUMMY_RESERVED 32'hffffffff
