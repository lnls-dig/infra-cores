package wb_acq_core_regs_consts_pkg is
  constant ADDR_ACQ_CORE_CTL : Natural := 16#0#;
  constant ACQ_CORE_CTL_FSM_START_ACQ_OFFSET : Natural := 0;
  constant ACQ_CORE_CTL_FSM_STOP_ACQ_OFFSET : Natural := 1;
  constant ACQ_CORE_CTL_RESERVED1_OFFSET : Natural := 2;
  constant ACQ_CORE_CTL_FSM_ACQ_NOW_OFFSET : Natural := 16;
  constant ACQ_CORE_CTL_RESERVED2_OFFSET : Natural := 17;
  constant ADDR_ACQ_CORE_STA : Natural := 16#4#;
  constant ACQ_CORE_STA_FSM_STATE_OFFSET : Natural := 0;
  constant ACQ_CORE_STA_FSM_ACQ_DONE_OFFSET : Natural := 3;
  constant ACQ_CORE_STA_FIFO_WE_OFFSET : Natural := 4;
  constant ACQ_CORE_STA_FIFO_RE_OFFSET : Natural := 5;
  constant ACQ_CORE_STA_FIFO_FC_RD_EN_OFFSET : Natural := 6;
  constant ACQ_CORE_STA_FIFO_RD_EMPTY_OFFSET : Natural := 7;
  constant ACQ_CORE_STA_FC_TRANS_DONE_OFFSET : Natural := 8;
  constant ACQ_CORE_STA_FC_FULL_OFFSET : Natural := 9;
  constant ACQ_CORE_STA_FIFO_WR_FULL_OFFSET : Natural := 10;
  constant ACQ_CORE_STA_FIFO_FC_VALID_FWFT_OFFSET : Natural := 11;
  constant ACQ_CORE_STA_SOURCE_PL_DREQ_OFFSET : Natural := 12;
  constant ACQ_CORE_STA_SOURCE_PL_STALL_OFFSET : Natural := 13;
  constant ACQ_CORE_STA_RESERVED2_OFFSET : Natural := 14;
  constant ACQ_CORE_STA_DDR3_TRANS_DONE_OFFSET : Natural := 16;
  constant ACQ_CORE_STA_FIFO_WR_COUNT_OFFSET : Natural := 17;
  constant ADDR_ACQ_CORE_TRIG_CFG : Natural := 16#8#;
  constant ACQ_CORE_TRIG_CFG_HW_TRIG_SEL_OFFSET : Natural := 0;
  constant ACQ_CORE_TRIG_CFG_HW_TRIG_POL_OFFSET : Natural := 1;
  constant ACQ_CORE_TRIG_CFG_HW_TRIG_EN_OFFSET : Natural := 2;
  constant ACQ_CORE_TRIG_CFG_SW_TRIG_EN_OFFSET : Natural := 3;
  constant ACQ_CORE_TRIG_CFG_INT_TRIG_SEL_OFFSET : Natural := 4;
  constant ACQ_CORE_TRIG_CFG_RESERVED_OFFSET : Natural := 9;
  constant ADDR_ACQ_CORE_TRIG_DATA_CFG : Natural := 16#c#;
  constant ACQ_CORE_TRIG_DATA_CFG_THRES_FILT_OFFSET : Natural := 0;
  constant ACQ_CORE_TRIG_DATA_CFG_RESERVED_OFFSET : Natural := 8;
  constant ADDR_ACQ_CORE_TRIG_DATA_THRES : Natural := 16#10#;
  constant ADDR_ACQ_CORE_TRIG_DLY : Natural := 16#14#;
  constant ADDR_ACQ_CORE_SW_TRIG : Natural := 16#18#;
  constant ADDR_ACQ_CORE_SHOTS : Natural := 16#1c#;
  constant ACQ_CORE_SHOTS_NB_OFFSET : Natural := 0;
  constant ACQ_CORE_SHOTS_MULTISHOT_RAM_SIZE_IMPL_OFFSET : Natural := 16;
  constant ACQ_CORE_SHOTS_MULTISHOT_RAM_SIZE_OFFSET : Natural := 17;
  constant ADDR_ACQ_CORE_TRIG_POS : Natural := 16#20#;
  constant ADDR_ACQ_CORE_PRE_SAMPLES : Natural := 16#24#;
  constant ADDR_ACQ_CORE_POST_SAMPLES : Natural := 16#28#;
  constant ADDR_ACQ_CORE_SAMPLES_CNT : Natural := 16#2c#;
  constant ADDR_ACQ_CORE_DDR3_START_ADDR : Natural := 16#30#;
  constant ADDR_ACQ_CORE_DDR3_END_ADDR : Natural := 16#34#;
  constant ADDR_ACQ_CORE_ACQ_CHAN_CTL : Natural := 16#38#;
  constant ACQ_CORE_ACQ_CHAN_CTL_WHICH_OFFSET : Natural := 0;
  constant ACQ_CORE_ACQ_CHAN_CTL_RESERVED_OFFSET : Natural := 5;
  constant ACQ_CORE_ACQ_CHAN_CTL_DTRIG_WHICH_OFFSET : Natural := 8;
  constant ACQ_CORE_ACQ_CHAN_CTL_RESERVED1_OFFSET : Natural := 13;
  constant ACQ_CORE_ACQ_CHAN_CTL_NUM_CHAN_OFFSET : Natural := 16;
  constant ACQ_CORE_ACQ_CHAN_CTL_RESERVED2_OFFSET : Natural := 21;
  constant ADDR_ACQ_CORE_CH0_DESC : Natural := 16#3c#;
  constant ACQ_CORE_CH0_DESC_INT_WIDTH_OFFSET : Natural := 0;
  constant ACQ_CORE_CH0_DESC_NUM_COALESCE_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH0_ATOM_DESC : Natural := 16#40#;
  constant ACQ_CORE_CH0_ATOM_DESC_NUM_ATOMS_OFFSET : Natural := 0;
  constant ACQ_CORE_CH0_ATOM_DESC_ATOM_WIDTH_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH1_DESC : Natural := 16#44#;
  constant ACQ_CORE_CH1_DESC_INT_WIDTH_OFFSET : Natural := 0;
  constant ACQ_CORE_CH1_DESC_NUM_COALESCE_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH1_ATOM_DESC : Natural := 16#48#;
  constant ACQ_CORE_CH1_ATOM_DESC_NUM_ATOMS_OFFSET : Natural := 0;
  constant ACQ_CORE_CH1_ATOM_DESC_ATOM_WIDTH_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH2_DESC : Natural := 16#4c#;
  constant ACQ_CORE_CH2_DESC_INT_WIDTH_OFFSET : Natural := 0;
  constant ACQ_CORE_CH2_DESC_NUM_COALESCE_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH2_ATOM_DESC : Natural := 16#50#;
  constant ACQ_CORE_CH2_ATOM_DESC_NUM_ATOMS_OFFSET : Natural := 0;
  constant ACQ_CORE_CH2_ATOM_DESC_ATOM_WIDTH_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH3_DESC : Natural := 16#54#;
  constant ACQ_CORE_CH3_DESC_INT_WIDTH_OFFSET : Natural := 0;
  constant ACQ_CORE_CH3_DESC_NUM_COALESCE_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH3_ATOM_DESC : Natural := 16#58#;
  constant ACQ_CORE_CH3_ATOM_DESC_NUM_ATOMS_OFFSET : Natural := 0;
  constant ACQ_CORE_CH3_ATOM_DESC_ATOM_WIDTH_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH4_DESC : Natural := 16#5c#;
  constant ACQ_CORE_CH4_DESC_INT_WIDTH_OFFSET : Natural := 0;
  constant ACQ_CORE_CH4_DESC_NUM_COALESCE_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH4_ATOM_DESC : Natural := 16#60#;
  constant ACQ_CORE_CH4_ATOM_DESC_NUM_ATOMS_OFFSET : Natural := 0;
  constant ACQ_CORE_CH4_ATOM_DESC_ATOM_WIDTH_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH5_DESC : Natural := 16#64#;
  constant ACQ_CORE_CH5_DESC_INT_WIDTH_OFFSET : Natural := 0;
  constant ACQ_CORE_CH5_DESC_NUM_COALESCE_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH5_ATOM_DESC : Natural := 16#68#;
  constant ACQ_CORE_CH5_ATOM_DESC_NUM_ATOMS_OFFSET : Natural := 0;
  constant ACQ_CORE_CH5_ATOM_DESC_ATOM_WIDTH_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH6_DESC : Natural := 16#6c#;
  constant ACQ_CORE_CH6_DESC_INT_WIDTH_OFFSET : Natural := 0;
  constant ACQ_CORE_CH6_DESC_NUM_COALESCE_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH6_ATOM_DESC : Natural := 16#70#;
  constant ACQ_CORE_CH6_ATOM_DESC_NUM_ATOMS_OFFSET : Natural := 0;
  constant ACQ_CORE_CH6_ATOM_DESC_ATOM_WIDTH_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH7_DESC : Natural := 16#74#;
  constant ACQ_CORE_CH7_DESC_INT_WIDTH_OFFSET : Natural := 0;
  constant ACQ_CORE_CH7_DESC_NUM_COALESCE_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH7_ATOM_DESC : Natural := 16#78#;
  constant ACQ_CORE_CH7_ATOM_DESC_NUM_ATOMS_OFFSET : Natural := 0;
  constant ACQ_CORE_CH7_ATOM_DESC_ATOM_WIDTH_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH8_DESC : Natural := 16#7c#;
  constant ACQ_CORE_CH8_DESC_INT_WIDTH_OFFSET : Natural := 0;
  constant ACQ_CORE_CH8_DESC_NUM_COALESCE_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH8_ATOM_DESC : Natural := 16#80#;
  constant ACQ_CORE_CH8_ATOM_DESC_NUM_ATOMS_OFFSET : Natural := 0;
  constant ACQ_CORE_CH8_ATOM_DESC_ATOM_WIDTH_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH9_DESC : Natural := 16#84#;
  constant ACQ_CORE_CH9_DESC_INT_WIDTH_OFFSET : Natural := 0;
  constant ACQ_CORE_CH9_DESC_NUM_COALESCE_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH9_ATOM_DESC : Natural := 16#88#;
  constant ACQ_CORE_CH9_ATOM_DESC_NUM_ATOMS_OFFSET : Natural := 0;
  constant ACQ_CORE_CH9_ATOM_DESC_ATOM_WIDTH_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH10_DESC : Natural := 16#8c#;
  constant ACQ_CORE_CH10_DESC_INT_WIDTH_OFFSET : Natural := 0;
  constant ACQ_CORE_CH10_DESC_NUM_COALESCE_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH10_ATOM_DESC : Natural := 16#90#;
  constant ACQ_CORE_CH10_ATOM_DESC_NUM_ATOMS_OFFSET : Natural := 0;
  constant ACQ_CORE_CH10_ATOM_DESC_ATOM_WIDTH_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH11_DESC : Natural := 16#94#;
  constant ACQ_CORE_CH11_DESC_INT_WIDTH_OFFSET : Natural := 0;
  constant ACQ_CORE_CH11_DESC_NUM_COALESCE_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH11_ATOM_DESC : Natural := 16#98#;
  constant ACQ_CORE_CH11_ATOM_DESC_NUM_ATOMS_OFFSET : Natural := 0;
  constant ACQ_CORE_CH11_ATOM_DESC_ATOM_WIDTH_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH12_DESC : Natural := 16#9c#;
  constant ACQ_CORE_CH12_DESC_INT_WIDTH_OFFSET : Natural := 0;
  constant ACQ_CORE_CH12_DESC_NUM_COALESCE_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH12_ATOM_DESC : Natural := 16#a0#;
  constant ACQ_CORE_CH12_ATOM_DESC_NUM_ATOMS_OFFSET : Natural := 0;
  constant ACQ_CORE_CH12_ATOM_DESC_ATOM_WIDTH_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH13_DESC : Natural := 16#a4#;
  constant ACQ_CORE_CH13_DESC_INT_WIDTH_OFFSET : Natural := 0;
  constant ACQ_CORE_CH13_DESC_NUM_COALESCE_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH13_ATOM_DESC : Natural := 16#a8#;
  constant ACQ_CORE_CH13_ATOM_DESC_NUM_ATOMS_OFFSET : Natural := 0;
  constant ACQ_CORE_CH13_ATOM_DESC_ATOM_WIDTH_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH14_DESC : Natural := 16#ac#;
  constant ACQ_CORE_CH14_DESC_INT_WIDTH_OFFSET : Natural := 0;
  constant ACQ_CORE_CH14_DESC_NUM_COALESCE_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH14_ATOM_DESC : Natural := 16#b0#;
  constant ACQ_CORE_CH14_ATOM_DESC_NUM_ATOMS_OFFSET : Natural := 0;
  constant ACQ_CORE_CH14_ATOM_DESC_ATOM_WIDTH_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH15_DESC : Natural := 16#b4#;
  constant ACQ_CORE_CH15_DESC_INT_WIDTH_OFFSET : Natural := 0;
  constant ACQ_CORE_CH15_DESC_NUM_COALESCE_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH15_ATOM_DESC : Natural := 16#b8#;
  constant ACQ_CORE_CH15_ATOM_DESC_NUM_ATOMS_OFFSET : Natural := 0;
  constant ACQ_CORE_CH15_ATOM_DESC_ATOM_WIDTH_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH16_DESC : Natural := 16#bc#;
  constant ACQ_CORE_CH16_DESC_INT_WIDTH_OFFSET : Natural := 0;
  constant ACQ_CORE_CH16_DESC_NUM_COALESCE_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH16_ATOM_DESC : Natural := 16#c0#;
  constant ACQ_CORE_CH16_ATOM_DESC_NUM_ATOMS_OFFSET : Natural := 0;
  constant ACQ_CORE_CH16_ATOM_DESC_ATOM_WIDTH_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH17_DESC : Natural := 16#c4#;
  constant ACQ_CORE_CH17_DESC_INT_WIDTH_OFFSET : Natural := 0;
  constant ACQ_CORE_CH17_DESC_NUM_COALESCE_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH17_ATOM_DESC : Natural := 16#c8#;
  constant ACQ_CORE_CH17_ATOM_DESC_NUM_ATOMS_OFFSET : Natural := 0;
  constant ACQ_CORE_CH17_ATOM_DESC_ATOM_WIDTH_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH18_DESC : Natural := 16#cc#;
  constant ACQ_CORE_CH18_DESC_INT_WIDTH_OFFSET : Natural := 0;
  constant ACQ_CORE_CH18_DESC_NUM_COALESCE_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH18_ATOM_DESC : Natural := 16#d0#;
  constant ACQ_CORE_CH18_ATOM_DESC_NUM_ATOMS_OFFSET : Natural := 0;
  constant ACQ_CORE_CH18_ATOM_DESC_ATOM_WIDTH_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH19_DESC : Natural := 16#d4#;
  constant ACQ_CORE_CH19_DESC_INT_WIDTH_OFFSET : Natural := 0;
  constant ACQ_CORE_CH19_DESC_NUM_COALESCE_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH19_ATOM_DESC : Natural := 16#d8#;
  constant ACQ_CORE_CH19_ATOM_DESC_NUM_ATOMS_OFFSET : Natural := 0;
  constant ACQ_CORE_CH19_ATOM_DESC_ATOM_WIDTH_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH20_DESC : Natural := 16#dc#;
  constant ACQ_CORE_CH20_DESC_INT_WIDTH_OFFSET : Natural := 0;
  constant ACQ_CORE_CH20_DESC_NUM_COALESCE_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH20_ATOM_DESC : Natural := 16#e0#;
  constant ACQ_CORE_CH20_ATOM_DESC_NUM_ATOMS_OFFSET : Natural := 0;
  constant ACQ_CORE_CH20_ATOM_DESC_ATOM_WIDTH_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH21_DESC : Natural := 16#e4#;
  constant ACQ_CORE_CH21_DESC_INT_WIDTH_OFFSET : Natural := 0;
  constant ACQ_CORE_CH21_DESC_NUM_COALESCE_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH21_ATOM_DESC : Natural := 16#e8#;
  constant ACQ_CORE_CH21_ATOM_DESC_NUM_ATOMS_OFFSET : Natural := 0;
  constant ACQ_CORE_CH21_ATOM_DESC_ATOM_WIDTH_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH22_DESC : Natural := 16#ec#;
  constant ACQ_CORE_CH22_DESC_INT_WIDTH_OFFSET : Natural := 0;
  constant ACQ_CORE_CH22_DESC_NUM_COALESCE_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH22_ATOM_DESC : Natural := 16#f0#;
  constant ACQ_CORE_CH22_ATOM_DESC_NUM_ATOMS_OFFSET : Natural := 0;
  constant ACQ_CORE_CH22_ATOM_DESC_ATOM_WIDTH_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH23_DESC : Natural := 16#f4#;
  constant ACQ_CORE_CH23_DESC_INT_WIDTH_OFFSET : Natural := 0;
  constant ACQ_CORE_CH23_DESC_NUM_COALESCE_OFFSET : Natural := 16;
  constant ADDR_ACQ_CORE_CH23_ATOM_DESC : Natural := 16#f8#;
  constant ACQ_CORE_CH23_ATOM_DESC_NUM_ATOMS_OFFSET : Natural := 0;
  constant ACQ_CORE_CH23_ATOM_DESC_ATOM_WIDTH_OFFSET : Natural := 16;
end package wb_acq_core_regs_consts_pkg;
