library work;
use work.fmc_adc_pkg.all;
use work.textio_extended_pkg.all;

-- dummy package declaration to satisfy compilers
package ifc_generic_pkg is
end ifc_generic_pkg;
