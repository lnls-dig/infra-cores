library work;
use work.fmc_adc_pkg.all;
use work.textio_extended_pkg.all;
