package wb_evt_cnt_regs_consts_pkg is
  constant c_WB_EVT_CNT_REGS_SIZE : Natural := 8;
  constant c_WB_EVT_CNT_REGS_CTL_ADDR : Natural := 16#0#;
  constant c_WB_EVT_CNT_REGS_CTL_TRIG_ACT_OFFSET : Natural := 0;
  constant c_WB_EVT_CNT_REGS_CNT_SNAP_ADDR : Natural := 16#4#;
end package wb_evt_cnt_regs_consts_pkg;
