`define ADDR_WB_TRIG_IFACE_CH0_CTL     10'h0
`define WB_TRIG_IFACE_CH0_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH0_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH0_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH0_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH0_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH0_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH0_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH0_CTL_TRANSM_COUNT_RST 32'h00000008
`define WB_TRIG_IFACE_CH0_CTL_POL_OFFSET 4
`define WB_TRIG_IFACE_CH0_CTL_POL 32'h00000010
`define ADDR_WB_TRIG_IFACE_CH0_CFG     10'h4
`define WB_TRIG_IFACE_CH0_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH0_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH0_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH0_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH0_COUNT   10'h8
`define WB_TRIG_IFACE_CH0_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH0_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH0_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH0_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH0_CFG_TRANSM_DELAY_LEN 10'hc
`define ADDR_WB_TRIG_IFACE_CH0_CFG_RCV_DELAY_LEN 10'h10
`define ADDR_WB_TRIG_IFACE_CH0_CFG_TRANSM_PULSE_TRAIN 10'h14
`define WB_TRIG_IFACE_CH0_CFG_TRANSM_PULSE_TRAIN_NUM_OFFSET 0
`define WB_TRIG_IFACE_CH0_CFG_TRANSM_PULSE_TRAIN_NUM 32'h0000ffff
`define WB_TRIG_IFACE_CH0_CFG_TRANSM_PULSE_TRAIN_RESERVED_OFFSET 16
`define WB_TRIG_IFACE_CH0_CFG_TRANSM_PULSE_TRAIN_RESERVED 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH1_CTL     10'h18
`define WB_TRIG_IFACE_CH1_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH1_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH1_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH1_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH1_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH1_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH1_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH1_CTL_TRANSM_COUNT_RST 32'h00000008
`define WB_TRIG_IFACE_CH1_CTL_POL_OFFSET 4
`define WB_TRIG_IFACE_CH1_CTL_POL 32'h00000010
`define ADDR_WB_TRIG_IFACE_CH1_CFG     10'h1c
`define WB_TRIG_IFACE_CH1_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH1_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH1_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH1_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH1_COUNT   10'h20
`define WB_TRIG_IFACE_CH1_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH1_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH1_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH1_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH1_CFG_TRANSM_DELAY_LEN 10'h24
`define ADDR_WB_TRIG_IFACE_CH1_CFG_RCV_DELAY_LEN 10'h28
`define ADDR_WB_TRIG_IFACE_CH1_CFG_TRANSM_PULSE_TRAIN 10'h2c
`define WB_TRIG_IFACE_CH1_CFG_TRANSM_PULSE_TRAIN_NUM_OFFSET 0
`define WB_TRIG_IFACE_CH1_CFG_TRANSM_PULSE_TRAIN_NUM 32'h0000ffff
`define WB_TRIG_IFACE_CH1_CFG_TRANSM_PULSE_TRAIN_RESERVED_OFFSET 16
`define WB_TRIG_IFACE_CH1_CFG_TRANSM_PULSE_TRAIN_RESERVED 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH2_CTL     10'h30
`define WB_TRIG_IFACE_CH2_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH2_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH2_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH2_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH2_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH2_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH2_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH2_CTL_TRANSM_COUNT_RST 32'h00000008
`define WB_TRIG_IFACE_CH2_CTL_POL_OFFSET 4
`define WB_TRIG_IFACE_CH2_CTL_POL 32'h00000010
`define ADDR_WB_TRIG_IFACE_CH2_CFG     10'h34
`define WB_TRIG_IFACE_CH2_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH2_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH2_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH2_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH2_COUNT   10'h38
`define WB_TRIG_IFACE_CH2_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH2_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH2_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH2_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH2_CFG_TRANSM_DELAY_LEN 10'h3c
`define ADDR_WB_TRIG_IFACE_CH2_CFG_RCV_DELAY_LEN 10'h40
`define ADDR_WB_TRIG_IFACE_CH2_CFG_TRANSM_PULSE_TRAIN 10'h44
`define WB_TRIG_IFACE_CH2_CFG_TRANSM_PULSE_TRAIN_NUM_OFFSET 0
`define WB_TRIG_IFACE_CH2_CFG_TRANSM_PULSE_TRAIN_NUM 32'h0000ffff
`define WB_TRIG_IFACE_CH2_CFG_TRANSM_PULSE_TRAIN_RESERVED_OFFSET 16
`define WB_TRIG_IFACE_CH2_CFG_TRANSM_PULSE_TRAIN_RESERVED 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH3_CTL     10'h48
`define WB_TRIG_IFACE_CH3_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH3_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH3_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH3_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH3_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH3_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH3_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH3_CTL_TRANSM_COUNT_RST 32'h00000008
`define WB_TRIG_IFACE_CH3_CTL_POL_OFFSET 4
`define WB_TRIG_IFACE_CH3_CTL_POL 32'h00000010
`define ADDR_WB_TRIG_IFACE_CH3_CFG     10'h4c
`define WB_TRIG_IFACE_CH3_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH3_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH3_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH3_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH3_COUNT   10'h50
`define WB_TRIG_IFACE_CH3_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH3_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH3_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH3_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH3_CFG_TRANSM_DELAY_LEN 10'h54
`define ADDR_WB_TRIG_IFACE_CH3_CFG_RCV_DELAY_LEN 10'h58
`define ADDR_WB_TRIG_IFACE_CH3_CFG_TRANSM_PULSE_TRAIN 10'h5c
`define WB_TRIG_IFACE_CH3_CFG_TRANSM_PULSE_TRAIN_NUM_OFFSET 0
`define WB_TRIG_IFACE_CH3_CFG_TRANSM_PULSE_TRAIN_NUM 32'h0000ffff
`define WB_TRIG_IFACE_CH3_CFG_TRANSM_PULSE_TRAIN_RESERVED_OFFSET 16
`define WB_TRIG_IFACE_CH3_CFG_TRANSM_PULSE_TRAIN_RESERVED 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH4_CTL     10'h60
`define WB_TRIG_IFACE_CH4_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH4_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH4_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH4_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH4_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH4_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH4_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH4_CTL_TRANSM_COUNT_RST 32'h00000008
`define WB_TRIG_IFACE_CH4_CTL_POL_OFFSET 4
`define WB_TRIG_IFACE_CH4_CTL_POL 32'h00000010
`define ADDR_WB_TRIG_IFACE_CH4_CFG     10'h64
`define WB_TRIG_IFACE_CH4_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH4_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH4_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH4_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH4_COUNT   10'h68
`define WB_TRIG_IFACE_CH4_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH4_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH4_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH4_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH4_CFG_TRANSM_DELAY_LEN 10'h6c
`define ADDR_WB_TRIG_IFACE_CH4_CFG_RCV_DELAY_LEN 10'h70
`define ADDR_WB_TRIG_IFACE_CH4_CFG_TRANSM_PULSE_TRAIN 10'h74
`define WB_TRIG_IFACE_CH4_CFG_TRANSM_PULSE_TRAIN_NUM_OFFSET 0
`define WB_TRIG_IFACE_CH4_CFG_TRANSM_PULSE_TRAIN_NUM 32'h0000ffff
`define WB_TRIG_IFACE_CH4_CFG_TRANSM_PULSE_TRAIN_RESERVED_OFFSET 16
`define WB_TRIG_IFACE_CH4_CFG_TRANSM_PULSE_TRAIN_RESERVED 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH5_CTL     10'h78
`define WB_TRIG_IFACE_CH5_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH5_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH5_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH5_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH5_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH5_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH5_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH5_CTL_TRANSM_COUNT_RST 32'h00000008
`define WB_TRIG_IFACE_CH5_CTL_POL_OFFSET 4
`define WB_TRIG_IFACE_CH5_CTL_POL 32'h00000010
`define ADDR_WB_TRIG_IFACE_CH5_CFG     10'h7c
`define WB_TRIG_IFACE_CH5_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH5_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH5_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH5_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH5_COUNT   10'h80
`define WB_TRIG_IFACE_CH5_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH5_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH5_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH5_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH5_CFG_TRANSM_DELAY_LEN 10'h84
`define ADDR_WB_TRIG_IFACE_CH5_CFG_RCV_DELAY_LEN 10'h88
`define ADDR_WB_TRIG_IFACE_CH5_CFG_TRANSM_PULSE_TRAIN 10'h8c
`define WB_TRIG_IFACE_CH5_CFG_TRANSM_PULSE_TRAIN_NUM_OFFSET 0
`define WB_TRIG_IFACE_CH5_CFG_TRANSM_PULSE_TRAIN_NUM 32'h0000ffff
`define WB_TRIG_IFACE_CH5_CFG_TRANSM_PULSE_TRAIN_RESERVED_OFFSET 16
`define WB_TRIG_IFACE_CH5_CFG_TRANSM_PULSE_TRAIN_RESERVED 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH6_CTL     10'h90
`define WB_TRIG_IFACE_CH6_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH6_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH6_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH6_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH6_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH6_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH6_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH6_CTL_TRANSM_COUNT_RST 32'h00000008
`define WB_TRIG_IFACE_CH6_CTL_POL_OFFSET 4
`define WB_TRIG_IFACE_CH6_CTL_POL 32'h00000010
`define ADDR_WB_TRIG_IFACE_CH6_CFG     10'h94
`define WB_TRIG_IFACE_CH6_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH6_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH6_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH6_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH6_COUNT   10'h98
`define WB_TRIG_IFACE_CH6_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH6_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH6_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH6_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH6_CFG_TRANSM_DELAY_LEN 10'h9c
`define ADDR_WB_TRIG_IFACE_CH6_CFG_RCV_DELAY_LEN 10'ha0
`define ADDR_WB_TRIG_IFACE_CH6_CFG_TRANSM_PULSE_TRAIN 10'ha4
`define WB_TRIG_IFACE_CH6_CFG_TRANSM_PULSE_TRAIN_NUM_OFFSET 0
`define WB_TRIG_IFACE_CH6_CFG_TRANSM_PULSE_TRAIN_NUM 32'h0000ffff
`define WB_TRIG_IFACE_CH6_CFG_TRANSM_PULSE_TRAIN_RESERVED_OFFSET 16
`define WB_TRIG_IFACE_CH6_CFG_TRANSM_PULSE_TRAIN_RESERVED 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH7_CTL     10'ha8
`define WB_TRIG_IFACE_CH7_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH7_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH7_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH7_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH7_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH7_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH7_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH7_CTL_TRANSM_COUNT_RST 32'h00000008
`define WB_TRIG_IFACE_CH7_CTL_POL_OFFSET 4
`define WB_TRIG_IFACE_CH7_CTL_POL 32'h00000010
`define ADDR_WB_TRIG_IFACE_CH7_CFG     10'hac
`define WB_TRIG_IFACE_CH7_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH7_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH7_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH7_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH7_COUNT   10'hb0
`define WB_TRIG_IFACE_CH7_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH7_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH7_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH7_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH7_CFG_TRANSM_DELAY_LEN 10'hb4
`define ADDR_WB_TRIG_IFACE_CH7_CFG_RCV_DELAY_LEN 10'hb8
`define ADDR_WB_TRIG_IFACE_CH7_CFG_TRANSM_PULSE_TRAIN 10'hbc
`define WB_TRIG_IFACE_CH7_CFG_TRANSM_PULSE_TRAIN_NUM_OFFSET 0
`define WB_TRIG_IFACE_CH7_CFG_TRANSM_PULSE_TRAIN_NUM 32'h0000ffff
`define WB_TRIG_IFACE_CH7_CFG_TRANSM_PULSE_TRAIN_RESERVED_OFFSET 16
`define WB_TRIG_IFACE_CH7_CFG_TRANSM_PULSE_TRAIN_RESERVED 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH8_CTL     10'hc0
`define WB_TRIG_IFACE_CH8_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH8_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH8_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH8_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH8_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH8_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH8_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH8_CTL_TRANSM_COUNT_RST 32'h00000008
`define WB_TRIG_IFACE_CH8_CTL_POL_OFFSET 4
`define WB_TRIG_IFACE_CH8_CTL_POL 32'h00000010
`define ADDR_WB_TRIG_IFACE_CH8_CFG     10'hc4
`define WB_TRIG_IFACE_CH8_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH8_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH8_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH8_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH8_COUNT   10'hc8
`define WB_TRIG_IFACE_CH8_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH8_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH8_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH8_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH8_CFG_TRANSM_DELAY_LEN 10'hcc
`define ADDR_WB_TRIG_IFACE_CH8_CFG_RCV_DELAY_LEN 10'hd0
`define ADDR_WB_TRIG_IFACE_CH8_CFG_TRANSM_PULSE_TRAIN 10'hd4
`define WB_TRIG_IFACE_CH8_CFG_TRANSM_PULSE_TRAIN_NUM_OFFSET 0
`define WB_TRIG_IFACE_CH8_CFG_TRANSM_PULSE_TRAIN_NUM 32'h0000ffff
`define WB_TRIG_IFACE_CH8_CFG_TRANSM_PULSE_TRAIN_RESERVED_OFFSET 16
`define WB_TRIG_IFACE_CH8_CFG_TRANSM_PULSE_TRAIN_RESERVED 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH9_CTL     10'hd8
`define WB_TRIG_IFACE_CH9_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH9_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH9_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH9_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH9_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH9_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH9_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH9_CTL_TRANSM_COUNT_RST 32'h00000008
`define WB_TRIG_IFACE_CH9_CTL_POL_OFFSET 4
`define WB_TRIG_IFACE_CH9_CTL_POL 32'h00000010
`define ADDR_WB_TRIG_IFACE_CH9_CFG     10'hdc
`define WB_TRIG_IFACE_CH9_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH9_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH9_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH9_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH9_COUNT   10'he0
`define WB_TRIG_IFACE_CH9_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH9_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH9_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH9_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH9_CFG_TRANSM_DELAY_LEN 10'he4
`define ADDR_WB_TRIG_IFACE_CH9_CFG_RCV_DELAY_LEN 10'he8
`define ADDR_WB_TRIG_IFACE_CH9_CFG_TRANSM_PULSE_TRAIN 10'hec
`define WB_TRIG_IFACE_CH9_CFG_TRANSM_PULSE_TRAIN_NUM_OFFSET 0
`define WB_TRIG_IFACE_CH9_CFG_TRANSM_PULSE_TRAIN_NUM 32'h0000ffff
`define WB_TRIG_IFACE_CH9_CFG_TRANSM_PULSE_TRAIN_RESERVED_OFFSET 16
`define WB_TRIG_IFACE_CH9_CFG_TRANSM_PULSE_TRAIN_RESERVED 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH10_CTL    10'hf0
`define WB_TRIG_IFACE_CH10_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH10_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH10_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH10_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH10_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH10_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH10_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH10_CTL_TRANSM_COUNT_RST 32'h00000008
`define WB_TRIG_IFACE_CH10_CTL_POL_OFFSET 4
`define WB_TRIG_IFACE_CH10_CTL_POL 32'h00000010
`define ADDR_WB_TRIG_IFACE_CH10_CFG    10'hf4
`define WB_TRIG_IFACE_CH10_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH10_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH10_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH10_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH10_COUNT  10'hf8
`define WB_TRIG_IFACE_CH10_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH10_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH10_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH10_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH10_CFG_TRANSM_DELAY_LEN 10'hfc
`define ADDR_WB_TRIG_IFACE_CH10_CFG_RCV_DELAY_LEN 10'h100
`define ADDR_WB_TRIG_IFACE_CH10_CFG_TRANSM_PULSE_TRAIN 10'h104
`define WB_TRIG_IFACE_CH10_CFG_TRANSM_PULSE_TRAIN_NUM_OFFSET 0
`define WB_TRIG_IFACE_CH10_CFG_TRANSM_PULSE_TRAIN_NUM 32'h0000ffff
`define WB_TRIG_IFACE_CH10_CFG_TRANSM_PULSE_TRAIN_RESERVED_OFFSET 16
`define WB_TRIG_IFACE_CH10_CFG_TRANSM_PULSE_TRAIN_RESERVED 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH11_CTL    10'h108
`define WB_TRIG_IFACE_CH11_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH11_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH11_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH11_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH11_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH11_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH11_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH11_CTL_TRANSM_COUNT_RST 32'h00000008
`define WB_TRIG_IFACE_CH11_CTL_POL_OFFSET 4
`define WB_TRIG_IFACE_CH11_CTL_POL 32'h00000010
`define ADDR_WB_TRIG_IFACE_CH11_CFG    10'h10c
`define WB_TRIG_IFACE_CH11_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH11_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH11_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH11_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH11_COUNT  10'h110
`define WB_TRIG_IFACE_CH11_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH11_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH11_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH11_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH11_CFG_TRANSM_DELAY_LEN 10'h114
`define ADDR_WB_TRIG_IFACE_CH11_CFG_RCV_DELAY_LEN 10'h118
`define ADDR_WB_TRIG_IFACE_CH11_CFG_TRANSM_PULSE_TRAIN 10'h11c
`define WB_TRIG_IFACE_CH11_CFG_TRANSM_PULSE_TRAIN_NUM_OFFSET 0
`define WB_TRIG_IFACE_CH11_CFG_TRANSM_PULSE_TRAIN_NUM 32'h0000ffff
`define WB_TRIG_IFACE_CH11_CFG_TRANSM_PULSE_TRAIN_RESERVED_OFFSET 16
`define WB_TRIG_IFACE_CH11_CFG_TRANSM_PULSE_TRAIN_RESERVED 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH12_CTL    10'h120
`define WB_TRIG_IFACE_CH12_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH12_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH12_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH12_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH12_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH12_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH12_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH12_CTL_TRANSM_COUNT_RST 32'h00000008
`define WB_TRIG_IFACE_CH12_CTL_POL_OFFSET 4
`define WB_TRIG_IFACE_CH12_CTL_POL 32'h00000010
`define ADDR_WB_TRIG_IFACE_CH12_CFG    10'h124
`define WB_TRIG_IFACE_CH12_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH12_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH12_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH12_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH12_COUNT  10'h128
`define WB_TRIG_IFACE_CH12_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH12_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH12_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH12_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH12_CFG_TRANSM_DELAY_LEN 10'h12c
`define ADDR_WB_TRIG_IFACE_CH12_CFG_RCV_DELAY_LEN 10'h130
`define ADDR_WB_TRIG_IFACE_CH12_CFG_TRANSM_PULSE_TRAIN 10'h134
`define WB_TRIG_IFACE_CH12_CFG_TRANSM_PULSE_TRAIN_NUM_OFFSET 0
`define WB_TRIG_IFACE_CH12_CFG_TRANSM_PULSE_TRAIN_NUM 32'h0000ffff
`define WB_TRIG_IFACE_CH12_CFG_TRANSM_PULSE_TRAIN_RESERVED_OFFSET 16
`define WB_TRIG_IFACE_CH12_CFG_TRANSM_PULSE_TRAIN_RESERVED 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH13_CTL    10'h138
`define WB_TRIG_IFACE_CH13_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH13_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH13_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH13_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH13_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH13_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH13_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH13_CTL_TRANSM_COUNT_RST 32'h00000008
`define WB_TRIG_IFACE_CH13_CTL_POL_OFFSET 4
`define WB_TRIG_IFACE_CH13_CTL_POL 32'h00000010
`define ADDR_WB_TRIG_IFACE_CH13_CFG    10'h13c
`define WB_TRIG_IFACE_CH13_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH13_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH13_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH13_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH13_COUNT  10'h140
`define WB_TRIG_IFACE_CH13_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH13_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH13_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH13_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH13_CFG_TRANSM_DELAY_LEN 10'h144
`define ADDR_WB_TRIG_IFACE_CH13_CFG_RCV_DELAY_LEN 10'h148
`define ADDR_WB_TRIG_IFACE_CH13_CFG_TRANSM_PULSE_TRAIN 10'h14c
`define WB_TRIG_IFACE_CH13_CFG_TRANSM_PULSE_TRAIN_NUM_OFFSET 0
`define WB_TRIG_IFACE_CH13_CFG_TRANSM_PULSE_TRAIN_NUM 32'h0000ffff
`define WB_TRIG_IFACE_CH13_CFG_TRANSM_PULSE_TRAIN_RESERVED_OFFSET 16
`define WB_TRIG_IFACE_CH13_CFG_TRANSM_PULSE_TRAIN_RESERVED 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH14_CTL    10'h150
`define WB_TRIG_IFACE_CH14_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH14_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH14_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH14_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH14_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH14_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH14_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH14_CTL_TRANSM_COUNT_RST 32'h00000008
`define WB_TRIG_IFACE_CH14_CTL_POL_OFFSET 4
`define WB_TRIG_IFACE_CH14_CTL_POL 32'h00000010
`define ADDR_WB_TRIG_IFACE_CH14_CFG    10'h154
`define WB_TRIG_IFACE_CH14_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH14_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH14_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH14_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH14_COUNT  10'h158
`define WB_TRIG_IFACE_CH14_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH14_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH14_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH14_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH14_CFG_TRANSM_DELAY_LEN 10'h15c
`define ADDR_WB_TRIG_IFACE_CH14_CFG_RCV_DELAY_LEN 10'h160
`define ADDR_WB_TRIG_IFACE_CH14_CFG_TRANSM_PULSE_TRAIN 10'h164
`define WB_TRIG_IFACE_CH14_CFG_TRANSM_PULSE_TRAIN_NUM_OFFSET 0
`define WB_TRIG_IFACE_CH14_CFG_TRANSM_PULSE_TRAIN_NUM 32'h0000ffff
`define WB_TRIG_IFACE_CH14_CFG_TRANSM_PULSE_TRAIN_RESERVED_OFFSET 16
`define WB_TRIG_IFACE_CH14_CFG_TRANSM_PULSE_TRAIN_RESERVED 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH15_CTL    10'h168
`define WB_TRIG_IFACE_CH15_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH15_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH15_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH15_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH15_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH15_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH15_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH15_CTL_TRANSM_COUNT_RST 32'h00000008
`define WB_TRIG_IFACE_CH15_CTL_POL_OFFSET 4
`define WB_TRIG_IFACE_CH15_CTL_POL 32'h00000010
`define ADDR_WB_TRIG_IFACE_CH15_CFG    10'h16c
`define WB_TRIG_IFACE_CH15_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH15_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH15_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH15_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH15_COUNT  10'h170
`define WB_TRIG_IFACE_CH15_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH15_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH15_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH15_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH15_CFG_TRANSM_DELAY_LEN 10'h174
`define ADDR_WB_TRIG_IFACE_CH15_CFG_RCV_DELAY_LEN 10'h178
`define ADDR_WB_TRIG_IFACE_CH15_CFG_TRANSM_PULSE_TRAIN 10'h17c
`define WB_TRIG_IFACE_CH15_CFG_TRANSM_PULSE_TRAIN_NUM_OFFSET 0
`define WB_TRIG_IFACE_CH15_CFG_TRANSM_PULSE_TRAIN_NUM 32'h0000ffff
`define WB_TRIG_IFACE_CH15_CFG_TRANSM_PULSE_TRAIN_RESERVED_OFFSET 16
`define WB_TRIG_IFACE_CH15_CFG_TRANSM_PULSE_TRAIN_RESERVED 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH16_CTL    10'h180
`define WB_TRIG_IFACE_CH16_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH16_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH16_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH16_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH16_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH16_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH16_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH16_CTL_TRANSM_COUNT_RST 32'h00000008
`define WB_TRIG_IFACE_CH16_CTL_POL_OFFSET 4
`define WB_TRIG_IFACE_CH16_CTL_POL 32'h00000010
`define ADDR_WB_TRIG_IFACE_CH16_CFG    10'h184
`define WB_TRIG_IFACE_CH16_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH16_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH16_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH16_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH16_COUNT  10'h188
`define WB_TRIG_IFACE_CH16_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH16_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH16_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH16_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH16_CFG_TRANSM_DELAY_LEN 10'h18c
`define ADDR_WB_TRIG_IFACE_CH16_CFG_RCV_DELAY_LEN 10'h190
`define ADDR_WB_TRIG_IFACE_CH16_CFG_TRANSM_PULSE_TRAIN 10'h194
`define WB_TRIG_IFACE_CH16_CFG_TRANSM_PULSE_TRAIN_NUM_OFFSET 0
`define WB_TRIG_IFACE_CH16_CFG_TRANSM_PULSE_TRAIN_NUM 32'h0000ffff
`define WB_TRIG_IFACE_CH16_CFG_TRANSM_PULSE_TRAIN_RESERVED_OFFSET 16
`define WB_TRIG_IFACE_CH16_CFG_TRANSM_PULSE_TRAIN_RESERVED 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH17_CTL    10'h198
`define WB_TRIG_IFACE_CH17_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH17_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH17_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH17_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH17_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH17_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH17_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH17_CTL_TRANSM_COUNT_RST 32'h00000008
`define WB_TRIG_IFACE_CH17_CTL_POL_OFFSET 4
`define WB_TRIG_IFACE_CH17_CTL_POL 32'h00000010
`define ADDR_WB_TRIG_IFACE_CH17_CFG    10'h19c
`define WB_TRIG_IFACE_CH17_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH17_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH17_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH17_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH17_COUNT  10'h1a0
`define WB_TRIG_IFACE_CH17_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH17_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH17_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH17_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH17_CFG_TRANSM_DELAY_LEN 10'h1a4
`define ADDR_WB_TRIG_IFACE_CH17_CFG_RCV_DELAY_LEN 10'h1a8
`define ADDR_WB_TRIG_IFACE_CH17_CFG_TRANSM_PULSE_TRAIN 10'h1ac
`define WB_TRIG_IFACE_CH17_CFG_TRANSM_PULSE_TRAIN_NUM_OFFSET 0
`define WB_TRIG_IFACE_CH17_CFG_TRANSM_PULSE_TRAIN_NUM 32'h0000ffff
`define WB_TRIG_IFACE_CH17_CFG_TRANSM_PULSE_TRAIN_RESERVED_OFFSET 16
`define WB_TRIG_IFACE_CH17_CFG_TRANSM_PULSE_TRAIN_RESERVED 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH18_CTL    10'h1b0
`define WB_TRIG_IFACE_CH18_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH18_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH18_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH18_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH18_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH18_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH18_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH18_CTL_TRANSM_COUNT_RST 32'h00000008
`define WB_TRIG_IFACE_CH18_CTL_POL_OFFSET 4
`define WB_TRIG_IFACE_CH18_CTL_POL 32'h00000010
`define ADDR_WB_TRIG_IFACE_CH18_CFG    10'h1b4
`define WB_TRIG_IFACE_CH18_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH18_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH18_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH18_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH18_COUNT  10'h1b8
`define WB_TRIG_IFACE_CH18_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH18_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH18_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH18_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH18_CFG_TRANSM_DELAY_LEN 10'h1bc
`define ADDR_WB_TRIG_IFACE_CH18_CFG_RCV_DELAY_LEN 10'h1c0
`define ADDR_WB_TRIG_IFACE_CH18_CFG_TRANSM_PULSE_TRAIN 10'h1c4
`define WB_TRIG_IFACE_CH18_CFG_TRANSM_PULSE_TRAIN_NUM_OFFSET 0
`define WB_TRIG_IFACE_CH18_CFG_TRANSM_PULSE_TRAIN_NUM 32'h0000ffff
`define WB_TRIG_IFACE_CH18_CFG_TRANSM_PULSE_TRAIN_RESERVED_OFFSET 16
`define WB_TRIG_IFACE_CH18_CFG_TRANSM_PULSE_TRAIN_RESERVED 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH19_CTL    10'h1c8
`define WB_TRIG_IFACE_CH19_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH19_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH19_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH19_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH19_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH19_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH19_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH19_CTL_TRANSM_COUNT_RST 32'h00000008
`define WB_TRIG_IFACE_CH19_CTL_POL_OFFSET 4
`define WB_TRIG_IFACE_CH19_CTL_POL 32'h00000010
`define ADDR_WB_TRIG_IFACE_CH19_CFG    10'h1cc
`define WB_TRIG_IFACE_CH19_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH19_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH19_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH19_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH19_COUNT  10'h1d0
`define WB_TRIG_IFACE_CH19_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH19_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH19_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH19_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH19_CFG_TRANSM_DELAY_LEN 10'h1d4
`define ADDR_WB_TRIG_IFACE_CH19_CFG_RCV_DELAY_LEN 10'h1d8
`define ADDR_WB_TRIG_IFACE_CH19_CFG_TRANSM_PULSE_TRAIN 10'h1dc
`define WB_TRIG_IFACE_CH19_CFG_TRANSM_PULSE_TRAIN_NUM_OFFSET 0
`define WB_TRIG_IFACE_CH19_CFG_TRANSM_PULSE_TRAIN_NUM 32'h0000ffff
`define WB_TRIG_IFACE_CH19_CFG_TRANSM_PULSE_TRAIN_RESERVED_OFFSET 16
`define WB_TRIG_IFACE_CH19_CFG_TRANSM_PULSE_TRAIN_RESERVED 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH20_CTL    10'h1e0
`define WB_TRIG_IFACE_CH20_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH20_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH20_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH20_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH20_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH20_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH20_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH20_CTL_TRANSM_COUNT_RST 32'h00000008
`define WB_TRIG_IFACE_CH20_CTL_POL_OFFSET 4
`define WB_TRIG_IFACE_CH20_CTL_POL 32'h00000010
`define ADDR_WB_TRIG_IFACE_CH20_CFG    10'h1e4
`define WB_TRIG_IFACE_CH20_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH20_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH20_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH20_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH20_COUNT  10'h1e8
`define WB_TRIG_IFACE_CH20_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH20_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH20_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH20_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH20_CFG_TRANSM_DELAY_LEN 10'h1ec
`define ADDR_WB_TRIG_IFACE_CH20_CFG_RCV_DELAY_LEN 10'h1f0
`define ADDR_WB_TRIG_IFACE_CH20_CFG_TRANSM_PULSE_TRAIN 10'h1f4
`define WB_TRIG_IFACE_CH20_CFG_TRANSM_PULSE_TRAIN_NUM_OFFSET 0
`define WB_TRIG_IFACE_CH20_CFG_TRANSM_PULSE_TRAIN_NUM 32'h0000ffff
`define WB_TRIG_IFACE_CH20_CFG_TRANSM_PULSE_TRAIN_RESERVED_OFFSET 16
`define WB_TRIG_IFACE_CH20_CFG_TRANSM_PULSE_TRAIN_RESERVED 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH21_CTL    10'h1f8
`define WB_TRIG_IFACE_CH21_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH21_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH21_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH21_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH21_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH21_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH21_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH21_CTL_TRANSM_COUNT_RST 32'h00000008
`define WB_TRIG_IFACE_CH21_CTL_POL_OFFSET 4
`define WB_TRIG_IFACE_CH21_CTL_POL 32'h00000010
`define ADDR_WB_TRIG_IFACE_CH21_CFG    10'h1fc
`define WB_TRIG_IFACE_CH21_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH21_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH21_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH21_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH21_COUNT  10'h200
`define WB_TRIG_IFACE_CH21_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH21_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH21_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH21_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH21_CFG_TRANSM_DELAY_LEN 10'h204
`define ADDR_WB_TRIG_IFACE_CH21_CFG_RCV_DELAY_LEN 10'h208
`define ADDR_WB_TRIG_IFACE_CH21_CFG_TRANSM_PULSE_TRAIN 10'h20c
`define WB_TRIG_IFACE_CH21_CFG_TRANSM_PULSE_TRAIN_NUM_OFFSET 0
`define WB_TRIG_IFACE_CH21_CFG_TRANSM_PULSE_TRAIN_NUM 32'h0000ffff
`define WB_TRIG_IFACE_CH21_CFG_TRANSM_PULSE_TRAIN_RESERVED_OFFSET 16
`define WB_TRIG_IFACE_CH21_CFG_TRANSM_PULSE_TRAIN_RESERVED 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH22_CTL    10'h210
`define WB_TRIG_IFACE_CH22_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH22_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH22_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH22_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH22_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH22_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH22_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH22_CTL_TRANSM_COUNT_RST 32'h00000008
`define WB_TRIG_IFACE_CH22_CTL_POL_OFFSET 4
`define WB_TRIG_IFACE_CH22_CTL_POL 32'h00000010
`define ADDR_WB_TRIG_IFACE_CH22_CFG    10'h214
`define WB_TRIG_IFACE_CH22_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH22_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH22_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH22_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH22_COUNT  10'h218
`define WB_TRIG_IFACE_CH22_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH22_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH22_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH22_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH22_CFG_TRANSM_DELAY_LEN 10'h21c
`define ADDR_WB_TRIG_IFACE_CH22_CFG_RCV_DELAY_LEN 10'h220
`define ADDR_WB_TRIG_IFACE_CH22_CFG_TRANSM_PULSE_TRAIN 10'h224
`define WB_TRIG_IFACE_CH22_CFG_TRANSM_PULSE_TRAIN_NUM_OFFSET 0
`define WB_TRIG_IFACE_CH22_CFG_TRANSM_PULSE_TRAIN_NUM 32'h0000ffff
`define WB_TRIG_IFACE_CH22_CFG_TRANSM_PULSE_TRAIN_RESERVED_OFFSET 16
`define WB_TRIG_IFACE_CH22_CFG_TRANSM_PULSE_TRAIN_RESERVED 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH23_CTL    10'h228
`define WB_TRIG_IFACE_CH23_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH23_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH23_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH23_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH23_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH23_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH23_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH23_CTL_TRANSM_COUNT_RST 32'h00000008
`define WB_TRIG_IFACE_CH23_CTL_POL_OFFSET 4
`define WB_TRIG_IFACE_CH23_CTL_POL 32'h00000010
`define ADDR_WB_TRIG_IFACE_CH23_CFG    10'h22c
`define WB_TRIG_IFACE_CH23_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH23_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH23_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH23_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH23_COUNT  10'h230
`define WB_TRIG_IFACE_CH23_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH23_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH23_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH23_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH23_CFG_TRANSM_DELAY_LEN 10'h234
`define ADDR_WB_TRIG_IFACE_CH23_CFG_RCV_DELAY_LEN 10'h238
`define ADDR_WB_TRIG_IFACE_CH23_CFG_TRANSM_PULSE_TRAIN 10'h23c
`define WB_TRIG_IFACE_CH23_CFG_TRANSM_PULSE_TRAIN_NUM_OFFSET 0
`define WB_TRIG_IFACE_CH23_CFG_TRANSM_PULSE_TRAIN_NUM 32'h0000ffff
`define WB_TRIG_IFACE_CH23_CFG_TRANSM_PULSE_TRAIN_RESERVED_OFFSET 16
`define WB_TRIG_IFACE_CH23_CFG_TRANSM_PULSE_TRAIN_RESERVED 32'hffff0000
